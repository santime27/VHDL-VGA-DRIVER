library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity message is
	Generic (   LW: INTEGER:=10;
				DW: INTEGER:=50;
				DL: INTEGER:=100;
				POSX: INTEGER:= 0;
			    POSY: INTEGER:= 0); 
   Port (       HCOUNT : in  STD_LOGIC_VECTOR (10 downto 0);
                VCOUNT : in  STD_LOGIC_VECTOR (10 downto 0);
                VALUE:   in  STD_LOGIC_VECTOR (3 downto 0);
                PAINT:   out  STD_LOGIC);
end message ;

architecture Behavioral of message is

    -- letras base de 10x20
    type char_bitmap is array (0 to 19) of STD_LOGIC_VECTOR(9 downto 0);
    
    constant CHAR_A: char_bitmap := (
        "000001111111111110000",
        "000111111111111111000",
        "011111111111111111111",
        "111111110000011111111",
        "111111110000011111111",
        "111111110000011111111",
        "111111111111111111111",
        "111111111111111111111",
        "111111110000011111111",
        "111111110000011111111"
    );

    constant CHAR_B: char_bitmap := (
    "111111111111111100000",
    "111111111111111110000",
    "111111111111111111111",
    "111111110000011111111",
    "111111111111111110000",
    "111111111111111100000",
    "111111111111111111000",
    "111111110000011111111",
    "111111111111111111111",
    "111111111111111111000"
    );

    constant CHAR_C: char_bitmap := (
        "000001111111111111111",
        "000111111111111111111",
        "011111111111111111111",
        "111111110000000000000",
        "111111110000000000000",
        "111111110000000000000",
        "111111110000000000000",
        "111111110000000000000",
        "011111111111111111111",
        "000111111111111111111"
    );

    constant CHAR_D: char_bitmap := (
        "111111111111111100000",
        "111111111111111111000",
        "111111111111111111111",
        "111111110000011111111",
        "111111110000011111111",
        "111111110000011111111",
        "111111110000011111111",
        "111111110000011111111",
        "111111111111111111111",
        "111111111111111111000"
    );

    constant CHAR_E: char_bitmap := (
        "111111111111111111111",
        "111111111111111111111",
        "111111111111111111111",
        "111111110000000000000",
        "111111111111111100000",
        "111111111111111100000",
        "111111111111111100000",
        "111111110000000000000",
        "111111111111111111111",
        "111111111111111111111"
    );

    constant CHAR_F: char_bitmap := (
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111000000000000",
        "11111111111111110000",
        "11111111111111110000",
        "11111111111111110000",
        "11111111000000000000",
        "11111111000000000000",
        "11111111000000000000"
    );

    constant CHAR_G: char_bitmap := (
        "00000111111111111111",
        "00011111111111111111",
        "01111111111111111111",
        "11111111000000000000",
        "11111111011111111111",
        "11111111011111111111",
        "11111111011111111111",
        "11111111000001111111",
        "01111111111111111111",
        "00011111111111111111"
    );

    constant CHAR_H: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111"
    );

    constant CHAR_I: char_bitmap := (
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111"
    );

    constant CHAR_J: char_bitmap := (
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "01111111111111111111",
        "00011111111111111100"
    );

    constant CHAR_K: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111111111111000",
        "11111111111111110000",
        "11111111111111111000",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111"
    );

    constant CHAR_L: char_bitmap := (
        "11111111000000000000",
        "11111111000000000000",
        "11111111000000000000",
        "11111111000000000000",
        "11111111000000000000",
        "11111111000000000000",
        "11111111000000000000",
        "11111111000000000000",
        "11111111111111111111",
        "11111111111111111111"
    );

    constant CHAR_M: char_bitmap := (
        "1111110000000011111",
        "11111111000001111111",
        "11111111110011111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111000101111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111"
    );

    constant CHAR_N: char_bitmap := (
        "1111110000001111111",
        "11111111000001111111",
        "11111111110001111111",
        "11111111111001111111",
        "11111111111111111111",
        "11111111001111111111",
        "11111111000111111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111"
    );

    constant CHAR_O: char_bitmap := (
        "00000111111111111000",
        "00011111111111111100",
        "01111111111111111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "01111111111111111111",
        "00011111111111111100"
    );

    constant CHAR_P: char_bitmap := (
        "11111111111111110000",
        "11111111111111111100",
        "11111111111111111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111111111111110",
        "11111111111111111000",
        "11111111000000000000",
        "11111111000000000000"
    );

    constant CHAR_Q: char_bitmap := (
        "00000111111111110000",
        "00011111111111111100",
        "01111111111111111110",
        "11111110000001111110",
        "11111110000001111110",
        "11111110000001111110",
        "11111110000001111110",
        "11111110000001111110",
        "01111111111111111111",
        "00011111111111111111"
    );

    constant CHAR_R: char_bitmap := (
        "11111111111111110000",
        "11111111111111111100",
        "11111111111111111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111111111111110",
        "11111111111111111110",
        "11111111000111111111",
        "11111111000001111111"
    );

    constant CHAR_S: char_bitmap := (
        "00000111111111111111",
        "00011111111111111111",
        "01111111111111111111",
        "11111111000000000000",
        "01111111111111110000",
        "00011111111111111000",
        "00000111111111111111",
        "00000000000001111111",
        "11111111111111111111",
        "11111111111111111100"
    );

    constant CHAR_T: char_bitmap := (
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "00000001111110000000",
        "00000001111110000000",
        "00000001111110000000",
        "00000001111110000000",
        "00000001111110000000",
        "00000001111110000000",
        "00000001111110000000"
    );

    constant CHAR_U: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "01111111111111111111",
        "00111111111111111100"
    );

    constant CHAR_V: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111111111111111",
        "11111111111111111100"
    );

    constant CHAR_W: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111001001111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111110111111111",
        "11111111000001111111"
    );

    constant CHAR_X: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "01111110000001111111",
        "00111111111111111000",
        "00001111111111110000",
        "00111111111111111000",
        "01111110000001111111",
        "11111111000001111111",
        "11111111000001111111"
    );

    constant CHAR_Y: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "01111110000001111111",
        "00111111111111111000",
        "00001111111111110000",
        "00000001111110000000",
        "00000001111110000000",
        "00000001111110000000",
        "00000001111110000000"
    );

    constant CHAR_Z: char_bitmap := (
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "00000001111111111111",
        "00000011111111111100",
        "00001111111111110000",
        "00011111111111100000",
        "00111111111111000000",
        "11111111111111111111",
        "11111111111111111111"
    );

    constant CHAR_1: char_bitmap := (
        "0000000000000111111",
        "0000000111111111111",
        "0011111111111111111",
        "1111111111111111111",
        "1111111111111111111",
        "1111111111111111111",
        "1111111111111111111",
        "1111111111111111111",
        "1111111111111111111",
        "1111111111111111111"
    );

    constant CHAR_2: char_bitmap := (
        "11111111111111110000",
        "11111111111111111100",
        "11111111111111111111",
        "00000000000001111111",
        "00000111111111111111",
        "00011111111111111000",
        "01111111111111110000",
        "11111111000000000000",
        "11111111111111111111",
        "11111111111111111111"
    );

    constant CHAR_3: char_bitmap := (
        "11111111111111110000",
        "11111111111111111000",
        "11111111111111111111",
        "00000000000001111111",
        "00000111111111111000",
        "00000111111111100000",
        "00000111111111111000",
        "00000000000001111111",
        "11111111111111111111",
        "11111111111111111100"
    );

    constant CHAR_4: char_bitmap := (
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111000001111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111"
    );

    constant CHAR_5: char_bitmap := (
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111000000000000",
        "11111111111111110000",
        "11111111111111111100",
        "11111111111111111111",
        "00000000000001111111",
        "11111111111111111111",
        "11111111111111111100"
    );

    constant CHAR_6: char_bitmap := (
        "0000011111111111111",
        "0001111111111111111",
        "0111111111111111111",
        "1111111100000000000",
        "1111111111111111000",
        "1111111111111111110",
        "1111111111111111111",
        "1111111100000111111",
        "0111111111111111111",
        "0001111111111111100"
    );

    constant CHAR_7: char_bitmap := (
        "11111111111111111111",
        "11111111111111111111",
        "11111111111111111111",
        "11111111000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111",
        "00000000000001111111"
    );

    constant CHAR_8: char_bitmap := (
        "00000111111111110000",
        "00011111111111111000",
        "01111111111111111111",
        "01111111000001111111",
        "00011111111111111110",
        "00000111111111110000",
        "00011111111111111110",
        "01111111000001111111",
        "01111111111111111111",
        "00011111111111111000"
    );

    constant CHAR_9: char_bitmap := (
        "00000111111111110000",
        "00011111111111111100",
        "01111111111111111111",
        "11111111000001111111",
        "01111111111111111111",
        "00011111111111111110",
        "00000111111111111111",
        "00000000000001111111",
        "11111111111111111111",
        "11111111111111111100"
);

	signal segments : STD_LOGIC_VECTOR (7 downto 0);
	signal xrectaneg : STD_LOGIC_VECTOR (10 downto 0);
	signal xrectaneg1 : STD_LOGIC_VECTOR (10 downto 0);
	signal xrectaneg2 : STD_LOGIC_VECTOR (10 downto 0);
	
	-- Constantes Geometricas Display
	-- Segmentos horizaontales
	constant SHX1 : INTEGER := POSX;
	constant SHX2 : INTEGER := POSX + DW;
	constant SHY1 : INTEGER := POSY;
	constant SHY2 : INTEGER := POSY + LW;
	constant SHY3 : INTEGER := POSY + DL/2 - LW/2;
	constant SHY4 : INTEGER := POSY + DL/2 + LW/2;
	constant SHY5 : INTEGER := POSY + DL - LW;
	constant SHY6 : INTEGER := POSY + DL;
	-- Segmentos Verticales
	constant SVY1 : INTEGER := POSY;
	constant SVY2 : INTEGER := POSY + DL/2 + LW/2;
	constant SVY3 : INTEGER := POSY + DL/2 - LW/2;
	constant SVY4 : INTEGER := POSY + DL;
	constant SVX1 : INTEGER := POSX;
	constant SVX2 : INTEGER := POSX + LW;
	constant SVX3 : INTEGER := POSX + DW - LW;
	constant SVX4 : INTEGER := POSX + DW;
begin

--	xrectapos <= ( ('0'&vcount(10 downto 1)) + (POSX+LW/2) - POSY/2);
--	xrectapos1 <= xrectapos - LW/2;
--	xrectapos2 <= xrectapos + LW/2;
	
	xrectaneg <= ( (POSX-LW/2+DW) + POSY/2 -('0'&vcount(10 downto 1)));
	xrectaneg1 <= xrectaneg - LW/2;
	xrectaneg2 <= xrectaneg + LW/2;
   with value select
	--          "abcdefgh"
   segments <= "11111101" when "0000",
					"11100000" when "0001",
					"11011010" when "0010",
					"11110010" when "0011",
					"01100110" when "0100",
					"10110110" when "0101",
					"10111110" when "0110",
					"11100000" when "0111",
					"11111110" when "1000",
					"11100110" when "1001",
					"11101110" when "1010",
					"00111100" when "1011",
					"10011100" when "1100",
					"01111100" when "1101",
					"10011110" when "1110",
					"10001110" when "1111",
					"00000000" when others;


	DIPLAY: process(segments,HCOUNT,VCOUNT,xrectaneg,xrectaneg2,xrectaneg1)
	begin
		-- segmento a
		if(segments(7)='1' and (HCOUNT>=SHX1)and(HCOUNT<=SHX2)and(VCOUNT>=SHY1)and(VCOUNT<=SHY2)) then
			PAINT <= '1';
		-- segmento g
		elsif (segments(1)='1' and (HCOUNT>=SHX1)and(HCOUNT<=SHX2)and(VCOUNT>=SHY3)and(VCOUNT<=SHY4)) then
			PAINT <= '1';
		-- segmento d
		elsif (segments(4)='1' and (HCOUNT>=SHX1)and(HCOUNT<=SHX2)and(VCOUNT>=SHY5)and(VCOUNT<=SHY6)) then
			PAINT <= '1';
		-- segmento b
		elsif (segments(6)='1' and (HCOUNT>=SVX3)and(HCOUNT<=SVX4)and(VCOUNT>=SVY1)and(VCOUNT<=SVY2)) then
			PAINT <= '1';
		-- segmento c
		elsif (segments(5)='1' and (HCOUNT>=SVX3)and(HCOUNT<=SVX4)and(VCOUNT>=SVY3)and(VCOUNT<=SVY4)) then
			PAINT <= '1';
		-- segmento f
		elsif (segments(2)='1' and (HCOUNT>=SVX1)and(HCOUNT<=SVX2)and(VCOUNT>=SVY1)and(VCOUNT<=SVY2)) then
			PAINT <= '1';
		-- segmento e
		elsif (segments(3)='1' and (HCOUNT>=SVX1)and(HCOUNT<=SVX2)and(VCOUNT>=SVY3)and(VCOUNT<=SVY4)) then
			PAINT <= '1';
		elsif ((segments(0)='1') and (HCOUNT>=xrectaneg1)and(HCOUNT<=xrectaneg2)and(VCOUNT>=SVY3)and(VCOUNT<=SVY4)) then
			PAINT <= '1';
		else
			PAINT <= '0';
		end if;
	end process;
end Behavioral;

